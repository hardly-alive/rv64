module regfile (
    input  logic        clk,
    input  logic        rst_n,

    // Read Ports
    input  logic [4:0]  rs1_addr_i,
    output logic [63:0] rs1_data_o,

    input  logic [4:0]  rs2_addr_i,
    output logic [63:0] rs2_data_o,

    // Write Port
    input  logic [4:0]  rd_addr_i,
    input  logic [63:0] rd_data_i,
    input  logic        rd_wen_i
);

    logic [63:0] regs [0:31];

    // ---------------------------------------------------------
    // WRITE LOGIC (Sequential)
    // ---------------------------------------------------------
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            for (int i=0; i<32; i++) regs[i] <= 64'b0;
        end else begin
            if (rd_wen_i && (rd_addr_i != 5'd0)) begin
                regs[rd_addr_i] <= rd_data_i;
            end
        end
    end

    // ---------------------------------------------------------
    // READ LOGIC (Combinational with Internal Forwarding)
    // ---------------------------------------------------------
    always_comb begin
        // Port 1
        if (rs1_addr_i == 5'd0) begin
            rs1_data_o = 64'b0;
        end else if ((rs1_addr_i == rd_addr_i) && rd_wen_i) begin
            // Forwarding: If writing to rs1 THIS CYCLE, output the new data immediately
            rs1_data_o = rd_data_i;
        end else begin
            rs1_data_o = regs[rs1_addr_i];
        end

        // Port 2
        if (rs2_addr_i == 5'd0) begin
            rs2_data_o = 64'b0;
        end else if ((rs2_addr_i == rd_addr_i) && rd_wen_i) begin
            rs2_data_o = rd_data_i;
        end else begin
            rs2_data_o = regs[rs2_addr_i];
        end
    end

endmodule