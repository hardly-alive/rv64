package riscv_pkg;

    // ------------------------------------
    // 1. Basic Parameters
    // ------------------------------------
    localparam int XLEN = 64;   // Data width
    localparam int ILEN = 32;   // Instruction width

    // ------------------------------------
    // 2. Opcodes (RV64I Base)
    // ------------------------------------
    typedef enum logic [6:0] {
        OP_LUI    = 7'b0110111,
        OP_AUIPC  = 7'b0010111,
        OP_JAL    = 7'b1101111,
        OP_JALR   = 7'b1100111,
        OP_BRANCH = 7'b1100011,
        OP_LOAD   = 7'b0000011,
        OP_STORE  = 7'b0100011,
        OP_IMM    = 7'b0010011, 
        OP_REG    = 7'b0110011,
        OP_SYSTEM = 7'b1110011 
    } opcode_t;

    // ------------------------------------
    // 3. ALU Operations
    // ------------------------------------
    typedef enum logic [3:0] {
        ALU_ADD,  ALU_SUB,
        ALU_SLL,  ALU_SLT,
        ALU_SLTU, ALU_XOR,
        ALU_SRL,  ALU_SRA,
        ALU_OR,   ALU_AND
    } alu_op_t;

endpackage